module fulladder (a,b);
